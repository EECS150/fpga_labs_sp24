module structural_adder (
    input [13:0] a,
    input [13:0] b,
    output [14:0] sum
);
    // TODO: Your implementation here.
    // TODO: Remove the assign statement below once you write your own RTL.
    assign sum = 15'd0;
endmodule
